`ifndef MACROS
`define MACROS

`define max(a, b) (((a) > (b)) ? (a) : (b))

`endif
